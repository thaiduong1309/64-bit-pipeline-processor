//Name1: Duong Bui
//Name2: Devin Stoen

module And(a, b, out);
					 
	input logic a, b;
	output logic out;
	
	and andgate2 (out, a, b);

endmodule