library verilog;
use verilog.vl_types.all;
entity mult_testbench is
end mult_testbench;
