library verilog;
use verilog.vl_types.all;
entity shifter_testbench is
end shifter_testbench;
