module STUR_REG(deout, writeData, d, dout);

	input logic [31:0][63:0] d;
	input logic [31:0]deout;
	input logic [63:0]writeData;
	output logic [31:0][63:0]dout;
	
	
	Stur_Reg[31:0][63:0];
	
	
	
	Stur_Reg[chooseREG][
	
	
	
	