library verilog;
use verilog.vl_types.all;
entity mux6432_1_testbench is
end mux6432_1_testbench;
